//Package file


`include "vm_seq_item.sv";
`include "vm_sequence.sv";
`include "vm_sequencer.sv";
`include "vm_monitor.sv";
`include "vm_driver.sv";
`include "vm_scoreboard.sv";
`include "vm_agent.sv";

`include "vm_env.sv";

`include "vm_test.sv";


